module Lessthan(in, out);
  input [31:0]in;
  output out;
 assign out = in[31];
endmodule