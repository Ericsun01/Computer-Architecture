module Overflow(input in1, input in2, output out);
	xor xorgate(out, in1, in2);
endmodule